library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
 

entity I_Memory is 
	port (addr: in std_logic_vector(15 downto 0); 
	
				data_read: out std_logic_vector(15 downto 0)
				);
end entity;

architecture Form of I_Memory is 
type ROMarray is array(100 downto 0) of std_logic_vector(7 downto 0);   -- defining a new type
signal ROM: ROMarray:=(0 =>"00010010",1 =>"10011000",
                       2 =>"00011111",3 =>"00110001",
                       4 =>"00010100",5 =>"10111010",
							  6 =>"00011000",7 =>"01100011",
							  8 =>"00010110",9 =>"10011100",
							  10 =>"00011011",11 =>"10111101",
							  12 =>"00011100",13 =>"01001110",
							  14 =>"00010100",15 =>"11001111",
							  16 =>"00101111",17 =>"00110001",
                       18 =>"00100100",19 =>"10111010",
							  20 =>"00101000",21 =>"01100011",
							  22 =>"00100110",23 =>"10011100",
							  24 =>"00101011",25 =>"10111101",
							  26 =>"00101100",27 =>"01001110",
							  28 =>"00001110",29 =>"10000001",
							  30 =>"00010011",31 =>"10000110",
                       32 =>"01011110",33 =>"10000100",
                       34 =>"01000010",35 =>"10000100",
							  36 =>"10001110",37 =>"11000001",
							  38 =>"10010011",39 =>"00000100",
							  40 =>"10101011",41 =>"11000100",
							  42 =>"11000100",43 =>"00000100",
                       44 =>"00010100",45 =>"11010100",
                       46 =>"01100100",47 =>"11010100",
							  48 =>"11000100",49 =>"00000100",
							  50 =>"11010101",51 =>"10000000",
							  others=>"00011000" );
signal d_read:std_logic_vector(15 downto 0):=(others=>'0');
begin
d_read(7 downto 0)<=ROM(to_integer(unsigned(addr))+1);
d_read(15 downto 8)<=ROM(to_integer(unsigned(addr)));	   	

data_read <= d_read;
	
	
	
end Form;